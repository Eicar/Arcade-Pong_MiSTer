/*
  MIT License

  Copyright (c) 2019 Richard Eng

  Permission is hereby granted, free of charge, to any person obtaining a copy
  of this software and associated documentation files (the "Software"), to deal
  in the Software without restriction, including without limitation the rights
  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
  copies of the Software, and to permit persons to whom the Software is
  furnished to do so, subject to the following conditions:

  The above copyright notice and this permission notice shall be included in all
  copies or substantial portions of the Software.

  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
  SOFTWARE.
*/

/*
  Pong - Vertical Sync Circuit
  ----------------------------
*/
`default_nettype none

module vsync
(
    input wire  mclk, vreset, v4, v8, v16,
    output wire vblank, _vblank, _vsync
);

srlatch f5cd(mclk, ~vreset, ~v16, vblank, _vblank);
assign _vsync = ~(vblank & v4 & ~v8);

/*
wire h5a_to_g5a;

wire _vblank_tmp;
ls02 f5c(vreset, vblank, _vblank_tmp);

reg _vblank_reg;
always @(posedge gclk) begin
  _vblank_reg <= _vblank_tmp;
end
assign _vblank = _vblank_reg;

wire vblank_tmp;
ls02 f5d(_vblank, v16, vblank_tmp);

reg vblank_reg;
always @(posedge gclk) begin
  vblank_reg <= vblank_tmp;
end
assign vblank = vblank_reg;

ls00 h5a(v8, v8, h5a_to_g5a);
ls10 g5a(vblank, v4, h5a_to_g5a, _vsync);
*/

endmodule
